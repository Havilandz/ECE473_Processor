// just the number 4

module four(
	output reg [31:0] four);
	
	always @* begin
		four <= 4;
	end
	
endmodule